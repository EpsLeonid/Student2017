package p;
	
	parameter SIZE_REG           = 8;

	parameter SIZE_DATA_OUT        = 16;

endpackage 