package parameters;
parameter reg_in = 7;
parameter reg_out = 15;
endpackage