package parmetry ;
    parameter sizeIn = 8 ;
    parameter sizeOut = 16;
endpackage 