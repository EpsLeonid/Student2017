package params;
	parameter INPUT_SIZE = 8;
	parameter STREAMS = 2;
	parameter OUTPUT_SIZE = 17;
endpackage
