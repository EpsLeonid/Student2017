package p_v5;  //параметры фильтра

	parameter k = 6;
	parameter l = 6;
	parameter M = 16;
endpackage