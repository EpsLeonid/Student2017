module D (

//------------------------------------------------------------
// Input Ports
//------------------------------------------------------------
	input  wire                                  clk,
	input  wire                                  d,
	

//------------------------------------------------------------
// Output Ports
//------------------------------------------------------------


	output  wire out);
	
	
	
	always @(posedge clk)
		begin
		out  <=d;
	end
endmodule