package v6_parametery_2;	 
	parameter k = 13;
	parameter l = 6;
	parameter m1 = 16;
	parameter m2 = 1;
	parameter size = k+l;
endpackage 