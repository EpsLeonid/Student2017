package v5_parameters;  //параметры фильтра

	parameter k = 6;
	parameter l = 6;
	parameter M = 16;
endpackage