import p::*; //параметризация
module R (

//------------------------------------------------------------
// входные порты
//------------------------------------------------------------
	input  wire                                  clk,
	input  reg [SIZE_REG - 1:0]                                 a,
	input  reg [SIZE_REG - 1:0]                                 b,
	input  reg [SIZE_REG - 1:0]                                 c,
	

//------------------------------------------------------------
// выходные порты
//------------------------------------------------------------

	output  reg [SIZE_DATA_OUT - 1:0]  DATA_OUT,
	output  reg [15:0]  s);
	
	//работа по клоку
	always @(posedge clk)
		begin
		s<=a*b;
		DATA_OUT  <=s+c;
	end
endmodule
	
