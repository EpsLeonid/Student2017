module D (

//------------------------------------------------------------
// входные порты
//------------------------------------------------------------
	input  wire                                  clk,
	input  wire                                  d,
	

//------------------------------------------------------------
// выходные порты
//------------------------------------------------------------


	output  wire out);
	
	
	//работа по клоку
	always @(posedge clk)
		begin
		out  <=d;
	end
endmodule
