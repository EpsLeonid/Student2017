package v4_parameters;	 
	parameter k = 9;
	parameter l = 5;
	parameter M = 6;
	parameter N = k + l;
endpackage 