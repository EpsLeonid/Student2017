module m (

//------------------------------------------------------------
// Input Ports
//------------------------------------------------------------
	input  wire                                  clk,
	input  wire                                  a,
	input  wire                                  b,


//------------------------------------------------------------
// Output Ports
//------------------------------------------------------------

	output  wire  c
);
	

	always @(posedge clk)
		begin
		c<=a*b;
	end
endmodule
