package settings;
parameter SIZE_REG_in = 8;
parameter SIZE_REG_out = 16;
endpackage 