package settings;
parameter SIZE_REG_1 = 8;
parameter SIZE_REG_2 = 16;
endpackage 