package param_P;

	parameter P=8;
	
endpackage 