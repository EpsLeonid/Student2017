package v8_parameters;  //параметры фильтра

	parameter k = 9;
	parameter l = 6;
	parameter M = 15;
endpackage