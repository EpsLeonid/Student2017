package V3_parameter;
	parameter l_3 = 5;
	parameter k_3 = 11;
	parameter m1 = 16;
	parameter m2 = 1;
endpackage
