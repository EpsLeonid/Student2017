package v1_filter_params;
	parameter M = 16;
	parameter k = 8;
	parameter l = 5;
endpackage
